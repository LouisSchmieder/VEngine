module opengl
