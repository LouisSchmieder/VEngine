module opengl

pub struct VAO {
}

pub fn new_vao() &VAO {
	return &VAO{}
}
