module mathf

pub struct Matrix {
mut:
	buffer [][]f32
}
