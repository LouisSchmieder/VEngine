module main

import backend
import backend.opengl

fn main() {
	mut backend := opengl.init_opengl()
}
